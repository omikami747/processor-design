module pc(
	  clk,
	  rst,
	  c_e,
	  adrs_in,
	  adrs_out,
	  en_pc
	  );
   input wire clk;
   input wire rst;
   input wire c_e;
   input wire [7:0] adrs_in;
   input wire 	    en_pc;
   
   output  wire [7:0] adrs_out;
   reg [7:0] 	    temp_adrs;
   
   always @(posedge clk or negedge rst)
     begin
	if(c_e & en_pc === 1'b0)
	  begin
	  end
	else if(rst === 1'b0)
	  begin
	     temp_adrs <= 8'b00000000;
	  end
	else
	  begin
	     temp_adrs <= adrs_in;
	  end
     end // always @ (posedge clk or negedge rst or negedge c_e)
   assign adrs_out = temp_adrs;
   
   
endmodule
