module toplevel(
		
		)
