module mux_a(
	     muxa,
	     acc,
	     pc,
	     a);
   
   input wire      muxa;
   input wire [7:0] acc;
   input wire [7:0]  pc;
   
   output reg [7:0] a;
   
   always @(*)
     begin
	if(muxa === 1'b0)
	  begin
	     a <= acc;
	  end
	else
	  begin
	     a <= pc;
	  end
     end // always @ (*)
   
endmodule // mux_a

